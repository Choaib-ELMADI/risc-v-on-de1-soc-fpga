module alu (ALUResult, Zero, ALUControl, SrcA, SrcB);
    output [31:0] ALUResult;
    output        Zero;
    input   [2:0] ALUControl;
    input  [31:0] SrcA, SrcB;

    // DO THE WORK HERE!

endmodule // alu
