module alu (
    input   [31:0] SrcA,
    input   [31:0] SrcB,
    input   [3:0]  aluc,
    output reg [31:0] Alu_out,
    output reg        zero,
    output reg        cout,
    output reg        overflow,
    output reg        sign
);
    // DO THE WORK HERE!

endmodule // alu
